///////////////////////////////////////////////////////////////////////////////////////////
// Tyler Anderson Wed, Apr 01, 2015 10:59:20 AM
//
// rs232_des.v
// "RS-232 Deserializer"
// A custom Verilog HDL module
//
// Deserialize RS-232 communication and handshake each character downstream
//   No flow control
//   No parity
//   1 stop bit
//
// Clock rate needs to be ~10x baud rate for this to really work
// 
///////////////////////////////////////////////////////////////////////////////////////////


module rs232_des
  (
   input 	    clk,     // clock frequency
   input 	    rst_n,   // active low reset
   input 	    rx,      // serial RS-232 data
   output reg [7:0] rx_data, // ascii data byte
   output reg 	    rx_req,  // request for downstream module to accept character
   input 	    rx_ack   // acknowledgement of acceptance from downstream
   );

`include "fncs.h"
   
   parameter P_CLK_FREQ_HZ = 100000000;
   parameter P_BAUD_RATE = 9600;

   // Goofy mark/space business
   wire 	    rx_n = !rx;
   
     
   // Finite state machine
   reg [1:0] 	    fsm;
   localparam
     S_IDLE  = 2'd0, // sit around waiting for a start bit
     S_START = 2'd1, // wait for the start bit to finish
     S_SHIFT = 2'd2, // shift in the serial data byte (little endian) and notify downstream when finished
     S_STOP  = 2'd3; // wait for the stop bit to finish
         
   // Synchronize rx into the clk domain and detect it's positive edgeOA
   wire 	    rx_n_s;
   wire 	    rx_n_s_pedge;
   sync SYNC0(.clk(clk), .rst_n(rst_n), .a(rx_n), .y(rx_n_s));
   posedge_detector PEDGE0(.clk(clk), .rst_n(rst_n), .a(rx_n_s), .y(rx_n_s_pedge));
   
   // Count to the center of each bit and latch on it
   localparam START_LATCH_CNT_MAX = P_CLK_FREQ_HZ/P_BAUD_RATE/2;
   localparam SHIFT_LATCH_CNT_MAX = P_CLK_FREQ_HZ/P_BAUD_RATE;
   localparam STOP_LATCH_CNT_MAX = P_CLK_FREQ_HZ/P_BAUD_RATE;
   localparam NBITS_LATCH_CNT = clogb2(SHIFT_LATCH_CNT_MAX);
   reg [NBITS_LATCH_CNT-1:0]  latch_cnt;

   // Count the 8 bits to be shifted in
   reg [2:0] 	    shift_cnt;

   // Handshake to downstream only if you get the stop bit (i.e., watch out for "break" condition.)
   // Note that downstream needs to be processing fast enough to keep up here
   always @(posedge clk or negedge rst_n )
     if( !rst_n ) rx_req <= 1'b0;
     else if( (fsm == S_STOP) && (latch_cnt == STOP_LATCH_CNT_MAX) && (rx_n_s == 1'b0) ) rx_req <= 1'b1;
     else if( rx_ack ) rx_req <= 1'b0;
     
   // Finite State Machine
   always @(posedge clk or negedge rst_n)
     if( !rst_n ) 
       begin
	  latch_cnt <= {NBITS_LATCH_CNT{1'b0}}; 
          shift_cnt <= 3'd0; 
	  rx_data <= 8'd0;
	  fsm <= S_IDLE;
       end
     
     else
       begin
	  case( fsm )
	    
	    S_IDLE:
	      begin
		 latch_cnt <= {NBITS_LATCH_CNT-1{1'b0}};
		 shift_cnt <= 3'd0;
		 if( rx_n_s_pedge )
		   fsm <= S_START;
	      end
		 
	    S_START: 
	      if( latch_cnt == START_LATCH_CNT_MAX )
		begin
		   latch_cnt <= {NBITS_LATCH_CNT-1{1'b0}}; 
	           fsm <= S_SHIFT; 
	        end
	      else 
                begin
		   latch_cnt <= latch_cnt + 1'b1;
		end
	    
	    S_SHIFT: 
	      if( (shift_cnt == 3'd7) && (latch_cnt == SHIFT_LATCH_CNT_MAX) )   
		begin
		   rx_data <= {rx_n_s,rx_data[7:1]}; // RS-232 is little endian
		   shift_cnt <= 3'b0;
		   latch_cnt <= {NBITS_LATCH_CNT-1{1'b0}}; 
		   fsm <= S_STOP;  
		end
	      else if( latch_cnt == SHIFT_LATCH_CNT_MAX )
		begin
		   rx_data <= {rx_n_s,rx_data[7:1]}; // RS-232 is little endian
		   shift_cnt <= shift_cnt + 1'b1;
		   latch_cnt <= {NBITS_LATCH_CNT-1{1'b0}};
		end
	      else
		begin
		   latch_cnt <= latch_cnt + 1'b1;
		end
	 
	    S_STOP:  
	      if( latch_cnt == STOP_LATCH_CNT_MAX  )   
		begin 
		   latch_cnt <= {NBITS_LATCH_CNT-1{1'b0}}; 
	           fsm <= S_IDLE;
	        end
	      else
		begin
		   latch_cnt <= latch_cnt + 1'b1;
		end

	    default: fsm <= S_IDLE;
	    
	  endcase // case ( fsm )
       end
   
endmodule // rs232_des

